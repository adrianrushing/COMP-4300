package delay_package is
    constant prop_delay : time := 5 ns;
end delay_package;